/*
 MIPS32 Core
 Designed by: danilo94
 This module have only one input and is used to contain all MIPS submodules 
*/
`include "ProgramCounter.v"


module mipsCore(input clk);















endmodule
