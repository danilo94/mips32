module mipsCore(input clk);















endmodule
