module Registers(input clk,
input [4:0] rs,
input [4:0] ra,
input [4:0] wr,
input [31:0] writeData,
input write,
output [31:0]readDatars,
output [31:0]readDatara);


reg [31:0] registers[0:31];

















endmodule
