controlUnity(
input [5:0] opcode,
output reg PCWrite,
output reg MemRead,
output reg MemWrite,
output reg MemtoReg,
output reg [1:0] PCSource,
output reg AluOp,
output reg AluScrcA,
output reg [2:0] AluSrcB,
output reg regWrite,
output reg regdst;
);













endmodule
